module test

pub fn my_print() {
	println('test')
}